
module instr_mem (
    input logic [31:0] addr,
    output logic [31:0] instruction
);

